`include "lib/defines.vh"
module WB(
    input wire clk,
    input wire rst,
    input wire [`StallBus-1:0] stall,
    input wire [`MEM_TO_WB_WD-1+64+1+2:0] mem_to_wb_bus,
    output wire [`WB_TO_RF_WD-1+64+1+2:0] wb_to_rf_bus,
    output wire [31:0] debug_wb_pc,
    output wire [3:0] debug_wb_rf_wen,
    output wire [4:0] debug_wb_rf_wnum,
    output wire [31:0] debug_wb_rf_wdata
    //

);

    reg [`MEM_TO_WB_WD-1+64+1+2:0] mem_to_wb_bus_r;

    always @ (posedge clk) begin
        if (rst) begin
            mem_to_wb_bus_r <= `MEM_TO_WB_WD+64+1+2'b0;
        end
        else if (stall[4]==`Stop && stall[5]==`NoStop) begin
            mem_to_wb_bus_r <= `MEM_TO_WB_WD+64+1+2'b0;
        end
        else if (stall[4]==`NoStop) begin
            mem_to_wb_bus_r <= mem_to_wb_bus;
        end
    end

    wire [31:0] wb_pc;
    wire rf_we;
    wire [4:0] rf_waddr;
    wire [31:0] rf_wdata;
    wire div_flag;
    wire [63:0] div_result;
    wire [1:0] mt_flag;
    
    assign {
        mt_flag,
        div_flag,         
        div_result,      
        wb_pc,
        rf_we,
        rf_waddr,
        rf_wdata
    } = mem_to_wb_bus_r;

//    assign wb_to_rf_bus = mem_to_wb_bus_r[`WB_TO_RF_WD-1:0];
    assign wb_to_rf_bus = {
        mt_flag,
        div_flag,         
        div_result,      
        rf_we,          //37
        rf_waddr,       //36:32
        rf_wdata        //31:0
    };

    assign debug_wb_pc = wb_pc;
    assign debug_wb_rf_wen = {4{rf_we}};
    assign debug_wb_rf_wnum = rf_waddr;
    assign debug_wb_rf_wdata = rf_wdata;

    
endmodule